library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity progmem IS
	port
	(
		address: in std_logic_vector (29 downto 0);
		clk: in std_logic  := '1';
		instruction_out: out std_logic_vector (31 downto 0)
	);
end progmem;


architecture behav of progmem is
	type rom_type is array (0 to 255) of std_logic_vector (31 downto 0);
	signal ROM : rom_type:=(
		-- Example program
		--x"00000000",
		--x"000027b7",
		--x"70f78513",
		--x"00100313",
		--x"00000293",
		--x"006283b3",
		--x"fea3dae3",
		--x"02702c23",
		--x"02602a23",
		--x"03402283",
	    --x"02702a23",
		--x"03402303",
		--x"fe5ff0ef",
		--x"00000001",
	 	--x"00000001",
		
		---------------------------------
		--Hazard Detection Unit
		--x"00000000",
		--x"03200293",
		--x"00400213",
		--x"04522823",
		--x"05022303",
		--x"05032303",
		--x"04600313",
		--x"05032383",
		--x"00040313",
		
		----------------------------------
		--x"00000000",
		--x"000022b7",
		--x"70f28293",
		--x"00001437",
		--x"d0540413",
		--x"04502823",
		--x"05002303",
		--x"408303b3",
		--x"05002303",
		--x"eb328493",
		---------------------------------
		--Rekursif
		x"00000000",
		x"40000113",
		x"090000ef",
		x"00050593",
		x"00a00893",

		x"00000013",
		x"fe010113",
		x"00112e23",
		x"00812c23",
		x"00912a23",		

		x"02010413",
		x"fea42623",
		x"fec42783",
		x"00079663",
		x"00000793",

		x"0440006f",
		x"fec42703",
		x"00100793",
		x"00f71663",
		x"00100793",
		
		x"0300006f",
		x"fec42783",
		x"fff78793",
		x"00078513",
		x"fb9ff0ef",

		x"00050493",
		x"fec42783",
		x"ffe78793",
		x"00078513",
		x"fa5ff0ef",		

		x"00050793",
		x"00f487b3",
		x"00078513",
		x"01c12083",
		x"01812403",

		x"01412483",
		x"02010113",
		x"00008067",
		x"fe010113",
		x"00112e23",	
		
		x"00812c23",
		x"02010413",
		x"fe042623",
		x"01400513",--00c00513
		x"00000097",		

		x"f68080e7",
		x"fea42623",
	
		x"00000013",
		x"ffdff06f",
		-----------
		--LUI
		--x"00000000",
		--x"0270f3b7",
		
		-----------
		--AUIPC
		--x"00000000",
		--x"00005397",
		-----------

		--BEQ
		--x"00000000",
		--x"00500293",
		--x"00028c63",
		--x"00000c63",
		--------------
		--BNE
	--	x"00000000",
		--x"00500293",
		--x"00001c63",
		--x"00029c63",
		--------------
		--BLT
		--x"00000000",
		--x"00500293",
		--x"0002cc63",
		--x"00504c63",
		--------------
		--BGE
		--x"00000000",
	--	x"00500293",
		--x"00505c63",
		--x"0002dc63",
		----------------
		--BLTU
		--x"00000000",
		--x"fff00293",
		--x"00506c63",
		--x"0002ec63",
		--------------
		--BGEU
		--x"00000000",
		--x"fff00293",
		--x"0002fc63",
		--x"00507c63",
		--------------
		--LB
		--x"00000000",
		--x"fff00293",
		--x"00502823",
		--x"01000303",
		--------------
		--LH
		--x"00000000",
		--x"fff00293",
		--x"00502823",
		--x"01001303",
		--------------
		--LW
		--x"00000000",
		--x"fff00293",
		--x"00502823",
		--x"01002303",
		--------------
		--LBU
		--x"00000000",
	--	x"fff00293",
	--	x"00502823",
	--	x"01004303",
		--------------
		--LHU
		--x"00000000",
	--	x"fff00293",
	--	x"00502823",
	--	x"01005303",
		--------------
		--SB
		--x"00000000",
	--	x"fff00293",
	--	x"00500823",
		--------------
		--SH
		--x"00000000",
		--x"fff00293",
		--x"00501823",
		--------------
		--SW
		--x"00000000",
		--x"fff00293",
		--x"00502823",
		--------------
		--ADDI
		--x"00000000",
		--x"fff00293",
		--------------
		--SLTI
		--x"00000000",
		--x"00200313",
		--x"00032293",
		--x"00332293",
		--------------
		--SLTIU
		--x"00000000",
		--x"00200313",
		--x"00033293",
		--x"00333293",
		--------------
		--XORI
		--x"00000000",
		--x"fff00293",
		--x"01f2c313",
		--------------
		--ORI
		--x"00000000",
		--x"ffff02b7",
		--x"10128293",
		--x"01f2e313",
		--------------
		--ANDI
		--x"00000000",
	--	x"ffff02b7",
	--	x"10128293",
		--x"01f2f313",
		--------------
		--SLLI
		--x"00000000",
		--x"ffff0337",
		--x"00331393",
		--------------
		--SRLI
		--x"00000000",
		--x"ffff0337",
		--x"00335393",
		--------------
		--SRAI
		--x"00000000",
		--x"ffff0337",
		--x"40335393",
		--------------
		--ADD
		--x"00000000",
	--	x"000102b7",
	--	x"fff28293",
	--	x"0000b337",
	--	x"bcd30313",
		--x"006283b3",
		--------------
		--SUB
		--x"00000000",
	--	x"000102b7",
	--	x"fff28293",
	--	x"0000b337",
	--	x"bcd30313",
	--	x"406283b3",
		--------------
		--SLL
		--x"00000000",
	--	x"ffff0337",
	--	x"ffff03b7",
	--	x"00138393",
	--	x"00731433",
		--------------
		--SLT
		--x"00000000",
	--	x"ffff0337",
	--	x"ffff03b7",
	--	x"00138393",
	--	x"00732433",
	--	x"0063a433",
		--------------
		--SLTU
		--x"00000000",
	--	x"ffff0337",
	--	x"ffff03b7",
	--	x"00138393",
	--	x"0063b433",
	--	x"00733433",
		--------------
		--XOR
		--x"00000000",
	--	x"000102b7",
	--	x"fff28293",
	--	x"0000b337",
	--	x"bcd30313",
	--	x"0062c3b3",
		--------------
		--SRL
		--x"00000000",
	--	x"ffff0337",
	--	x"ffff03b7",
	--	x"00138393",
	--	x"00735433",
		--------------
		--SRA
		--x"00000000",
	--	x"ffff0337",
	--	x"ffff03b7",
	--	x"00138393",
	--	x"40735433",
		--------------
		--OR
		--x"00000000",
	--	x"000102b7",
	--	x"fff28293",
	--	x"0000b337",
	--	x"bcd30313",
	--	x"0062e3b3",
		--------------
		--AND
		--x"00000000",
	--	x"000102b7",
	--	x"fff28293",
	--	x"0000b337",
	--	x"bcd30313",
	--	x"0062f3b3",
		
		--JAL
		--x"00000000",
	--	x"030000ef",
		------------
		--JALR
		--x"00000000",
	--	x"00c00293",
	--	x"00c28367",
		-------------
		others => x"00000000"
	);
begin
	instruction_out <= ROM(to_integer(unsigned(address)));
end behav;